
interface d_if ();

	logic clk;
	logic reset;
	logic d;
	logic q;
	logic qb;
	
endinterface : d_if

